    Mac OS X            	   2   �                                           ATTR         �   X                  �     com.apple.lastuseddate#PS       �   H  com.apple.macl   �2f    6�E     zu�ߊG��C�                                                      