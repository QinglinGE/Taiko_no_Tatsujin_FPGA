`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 05/01/2024 01:51:59 AM
// Design Name: 
// Module Name: music_rom
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module music_rom( 
    input logic[9:0]addr,
    output logic[7:0]data);
    parameter [0:280][7:0] ROM = {
    8'b01000000,
    //1
    8'b01111001,//1`
    8'b01111001,//1`
    //2
    8'b01111001,//1`
    8'b01111011,//3`
    //3
    8'b01111110,//6`
    8'b01111110,//6`
    //4
    8'b01111110,//6`
    8'b01111101,//5`
    //5
    8'b01111011,//3`
    8'b01111011,//3`
    //6
    8'b01111011,//3`
    8'b01111011,//3`
    //7
    8'b01110111,//7`,
    8'b01110111,//7`
    //8
    8'b01110111,//7`
    8'b01110110,//6`
    //9
    8'b01111001,//1`
    8'b01111001,//1`
    //10
    8'b01111001,//1`
    8'b01111011,//3`
    //11
    8'b01111110,//6`
    8'b01111110,//6`
    //12
    8'b01111110,//6`
    8'b01111101,//5`
    //13
    8'b01111011,//3`
    8'b01111011,//3`
    //14
    8'b01111011,//3`
    8'b01111011,//3`
    //15
    8'b01110111,//7
    8'b01110111,//7
    //16*4+1
    8'b01110111,//7
    8'b01110110,//6
    //72
    8'b01100000,
    8'b00111001,//1`
    8'b00111001,//1`
    8'b00110110,//6
    8'b00111001,//1`
    8'b00110110,//6
    8'b00111001,//1`
    8'b00111010,//2`
    //77
    8'b01111011,//3`
    8'b00111001,//1`
    8'b00111001,//1`
    8'b00110101,//5
    8'b01011011,//3` fudian
    //83
    8'b01100000,
    8'b01100000,
    8'b00100000,
    8'b00111001,//1`
    8'b00111001,//1`
    8'b00111001,//1`
    //88
    8'b01010111,//7 fudian
    8'b00110111,//7
    8'b00110110,//6
    8'b00110110,//6
    8'b01111001,//1`
    
    8'b01100000,
    8'b00111001,//1`
    8'b00111001,//1`
    8'b00110110,//6
    8'b00111001,//1`
    8'b00110110,//6
    8'b00111001,//1`
    8'b00111010,//2`
    //77
    8'b01111011,//3`
    8'b00111001,//1`
    8'b00111001,//1`
    8'b00111101,//5
    8'b01011011,//3` fudian
    //83
    8'b01100000,
    8'b01100000,
    8'b00100000,
    8'b00111001,//1`
    8'b00111001,//1`
    8'b01011010,//2`
    //88
    8'b01110000,
    8'b00110000,
    8'b00111011,//3`
    8'b00111011,//3`
    8'b00111011,//3`
    //
    8'b01111011,//3`
    8'b01110001,//1
    8'b01110001,//1
    8'b01110011,//3
    //
    8'b01110110,//6
    8'b01110110,//6
    8'b00110110,//6
    8'b00111011,//3`
    8'b00111011,//3`
    8'b00111011,//3`
    //
    8'b01111011,//3`
    8'b01111011,//3`
    8'b01111011,//3`
    8'b01111011,//3`
    //
    8'b01110111,//7
    8'b01110111,//7
    8'b00110111,//7
    8'b00111011,//3`
    8'b00111011,//3`
    8'b00111011,//3`
    //
    8'b01111011,//3'
    8'b01111001,//1`
    8'b00111001,//1`
    8'b00111010,//2`
    8'b00111010,//2`
    8'b00011010,//2`
    8'b00011011,//3`
    //
    8'b00111010,//2'
    8'b00111001,//1`
    8'b01111001,//1`
    8'b00110110,//6
    8'b00111011,//3`
    8'b00111011,//3`
    8'b00111011,//3`
    //
    8'b01111011,//3`
    8'b01111011,//3`
    8'b00111011,//3`
    8'b00111001,//1`
    8'b00111001,//1`
    8'b00011001,//1`
    8'b00011010,//2`
    //
    8'b00110111,//7
    8'b00110111,//7
    8'b00110111,//7
    8'b00111001,//1`
    8'b01111001,//1`
    8'b01100000,//
    //
    8'b00100000,//
    8'b00111011,//3`
    8'b00111011,//3`
    8'b00111011,//3`
    8'b11111011,//3`
    8'b01100000,//
    8'b00100000,//
    8'b00111001,//1`
    //
    8'b00110110,//6
    8'b11110101,//5
    8'b00111001,//1`
    8'b00111101,//5'
    8'b00011101,//5'
    8'b00011011,//3'
    //
    8'b11111011,//3'
    8'b00100000,//0'
    8'b00111001,//1`
    8'b00111101,//5'
    8'b00011101,//5'
    8'b00011010,//2`
    //
    8'b01111010,//2`
    8'b01100000,//
    8'b00100000,//0'
    8'b00111011,//3`
    8'b00111011,//3`
    8'b00111011,//3`
    //
    8'b11111011,//3`
    8'b00100000,//
    8'b00111001,//1`
    8'b00110110,//6
    8'b00010110,//6
    8'b00011100,//4'
    //
    8'b11111100,//4'
    8'b01100000,//0
    8'b00100000,//0
    8'b00111101,//5'
    //
    8'b00111011,//3`
    8'b00111101,//5'
    8'b00111011,//3`
    8'b00111101,//5'
    8'b00111011,//3`
    8'b00111101,//5'
    8'b00111011,//3`
    8'b00011011,//3`
    8'b01011100,//4'
    //
    8'b01110111,//7
    8'b01111100,//4'
    8'b01111011,//3'
    8'b01111001,//1`
    8'b01111001,//1`
    //2
    8'b01111001,//1`
    8'b01111011,//3`
    //3
    8'b01111110,//6`
    8'b01111110,//6`
    //4
    8'b01111110,//6`
    8'b01111101,//5`
    //5
    8'b01111011,//3`
    8'b01111011,//3`
    //6
    8'b01111011,//3`
    8'b01111011,//3`
    //7
    8'b01110111,//7`,
    8'b01110111,//7`
    //8
    8'b01110111,//7`
    8'b01110110,//6`
    8'b01111001,//1`
    8'b01111001,//1`
    //2
    8'b01111001,//1`
    8'b01111011,//3`
    //3
    8'b01111110,//6`
    8'b01111110,//6`
    //4
    8'b01111110,//6`
    8'b01111101,//5`
    //5
    8'b01111011,//3`
    8'b01111011,//3`
    //6
    8'b01111011,//3`
    8'b01111011,//3`
    //7
    8'b01110111,//7`,
    8'b01110111,//7`
    //8
    8'b01110111,//7`
    8'b01110110//6`
    
//test   
//      8'b10000000,
//      8'b10000001,
//      8'b10000010,
//      8'b10000011,
      
//      8'b10000100,
//      8'b10000101,
//      8'b10000110,
//      8'b10000111,
      
//      8'b00001000,
//      8'b00001001,
//      8'b00001010,
//      8'b00001011,
      
//      8'b01001100,
//      8'b01001101,
//      8'b01001110,
//      8'b01001111,
      
//      8'b01000000,
//      8'b01000001,
//      8'b01000010,
//      8'b01000011,
      
//      8'b01000100,
//      8'b01000101
  
    };
    assign data = ROM[addr];
endmodule
